module main;
	initial begin
	$display("hello from verilog");
	$finish;
	end
endmodule